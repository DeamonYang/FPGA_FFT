library verilog;
use verilog.vl_types.all;
entity fft_tb is
end fft_tb;
